module and_module (
    input a,
    input b,
    output c
);//{
    assign c = a & b; // And of two inputs
endmodule //}
